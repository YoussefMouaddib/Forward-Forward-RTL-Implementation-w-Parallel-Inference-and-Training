// tb_top.sv
// Testbench for neural_network_top.sv
// Simulates complete Forward-Forward training loop.
//
// RESPONSIBILITIES:
//   1. Load MNIST images and labels from .mem files
//   2. Instantiate DUT (neural_network_top)
//   3. Initialize weight BRAMs with Python-exported initial weights
//   4. Drive clock and reset
//   5. Monitor training progress via $display
//   6. Checkpoint weights periodically — dump to .mem files
//   7. Log goodness values and sample count for learning curve
//   8. Verify done signal and report final state
//
// VERIFICATION STRATEGY:
//   Primary: weight values change during training (learning happening)
//   Secondary: goodness separation visible in log
//   Against: Python golden reference output
//
// MEM FILE FORMAT:
//   All Q16.16, 32-bit hex, one value per line
//   Generated by ff_reference.py export_weights_to_mem()
//
// SIMULATION TIME:
//   At 100MHz, one sample takes roughly 1.2M cycles
//   7000 samples = 8.4B cycles — too slow for full RTL sim
//   Use NUM_SAMPLES=100 for functional verification
//   Scale up once verified correct

`timescale 1ns/1ps

module tb_top;

    // ─────────────────────────────────────────────
    // PARAMETERS
    // Match DUT parameters exactly
    // Use small sample count for simulation speed
    // ─────────────────────────────────────────────
    localparam L1_INPUT_SIZE  = 784;
    localparam L1_NUM_NEURONS = 256;
    localparam L2_INPUT_SIZE  = 256;
    localparam L2_NUM_NEURONS = 256;
    localparam DATA_WIDTH     = 32;
    localparam FRAC_BITS      = 16;
    localparam NUM_SAMPLES    = 100;   // small for sim — change to 7000 for full run
    localparam L1_DEPTH       = L1_NUM_NEURONS * L1_INPUT_SIZE;
    localparam L2_DEPTH       = L2_NUM_NEURONS * L2_INPUT_SIZE;

    // Checkpoint interval — dump weights every N samples
    localparam CHECKPOINT_INTERVAL = 10;

    // ─────────────────────────────────────────────
    // CLOCK AND RESET
    // ─────────────────────────────────────────────
    logic clk;
    logic rst_n;
    logic start;
    logic training_done;

    // 100MHz clock — 10ns period
    initial clk = 0;
    always #5 clk = ~clk;

    // ─────────────────────────────────────────────
    // SAMPLE AND LABEL MEMORIES
    // Loaded from Python-generated .mem files
    // Sized for NUM_SAMPLES images
    // ─────────────────────────────────────────────
    logic [0:(NUM_SAMPLES * L1_INPUT_SIZE)-1][DATA_WIDTH-1:0] sample_mem ;
    logic [0:NUM_SAMPLES-1][3:0]            label_mem  ;

    // DUT memory interface wires
    logic [$clog2(NUM_SAMPLES * L1_INPUT_SIZE)-1:0] sample_addr;
    logic        sample_en;
    logic [DATA_WIDTH-1:0] sample_rdata;
    logic [$clog2(NUM_SAMPLES)-1:0] label_addr;
    logic        label_en;
    logic [3:0]  label_rdata;

    // Memory read — synchronous to match DUT expectation
    always_ff @(posedge clk) begin
        if (sample_en)
            sample_rdata <= sample_mem[sample_addr];
        if (label_en)
            label_rdata <= label_mem[label_addr];
    end

    // ─────────────────────────────────────────────
    // DUT INSTANTIATION
    // ─────────────────────────────────────────────
    neural_network_top #(
        .L1_INPUT_SIZE  (L1_INPUT_SIZE),
        .L1_NUM_NEURONS (L1_NUM_NEURONS),
        .L2_INPUT_SIZE  (L2_INPUT_SIZE),
        .L2_NUM_NEURONS (L2_NUM_NEURONS),
        .DATA_WIDTH     (DATA_WIDTH),
        .FRAC_BITS      (FRAC_BITS),
        .NUM_SAMPLES    (NUM_SAMPLES)
    ) dut (
        .clk          (clk),
        .rst_n        (rst_n),
        .start        (start),
        .training_done(training_done),
        .sample_addr  (sample_addr),
        .sample_en    (sample_en),
        .sample_rdata (sample_rdata),
        .label_addr   (label_addr),
        .label_en     (label_en),
        .label_rdata  (label_rdata)
    );

    // ─────────────────────────────────────────────
    // WEIGHT INITIALIZATION
    // Load Python-exported initial weights into
    // DUT weight BRAMs using hierarchical references
    // This is testbench-only — not synthesizable
    // ─────────────────────────────────────────────
    task load_weights();
        $display("[TB] Loading initial weights from mem_files/...");
        $readmemh("C:/Users/youss/Documents/Forward-Forward-RTL-Implementation-w-Parallel-Inference-and-Training/mem_files/initial_layer1_w.mem", dut.l1_wbram.mem);
        $readmemh("C:/Users/youss/Documents/Forward-Forward-RTL-Implementation-w-Parallel-Inference-and-Training/mem_files/initial_layer2_w.mem", dut.l2_wbram.mem);
        $readmemh("C:/Users/youss/Documents/Forward-Forward-RTL-Implementation-w-Parallel-Inference-and-Training/mem_files/initial_layer1_b.mem", dut.l1_bias);
        $readmemh("C:/Users/youss/Documents/Forward-Forward-RTL-Implementation-w-Parallel-Inference-and-Training/mem_files/initial_layer2_b.mem", dut.l2_bias);
        $display("[TB] Weights loaded.");
    endtask

    // ─────────────────────────────────────────────
    // WEIGHT CHECKPOINT
    // Dump current weight BRAM contents to file
    // Call periodically to track learning
    // Compare against Python reference offline
    // ─────────────────────────────────────────────
    integer checkpoint_num;

    task dump_weights(input integer chk_num);
        string fname_l1, fname_l2;
        $sformat(fname_l1, "checkpoints/chk%0d_layer1_w.mem", chk_num);
        $sformat(fname_l2, "checkpoints/chk%0d_layer2_w.mem", chk_num);
        $writememh(fname_l1, dut.l1_wbram.mem);
        $writememh(fname_l2, dut.l2_wbram.mem);
        $display("[TB] Checkpoint %0d written at sample %0d",
                 chk_num, chk_num * CHECKPOINT_INTERVAL);
    endtask

    // ─────────────────────────────────────────────
    // GOODNESS MONITOR
    // Watches goodness values as they are produced
    // Logs to console and to file for plotting
    // ─────────────────────────────────────────────
    integer log_file;
    real    pos_goodness_f, neg_goodness_f;

    // Convert Q16.16 to real for display
    function real q_to_real(input logic signed [DATA_WIDTH-1:0] q);
        q_to_real = $itor($signed(q)) / 65536.0;
    endfunction

    // Monitor goodness_l2 done signal
    // When it fires, log current goodness values
    logic prev_goodness_l2_done;
    logic prev_goodness_l1_done;
    integer sample_count;
    logic   in_positive_pass;

    always_ff @(posedge clk) begin
        prev_goodness_l1_done <= dut.goodness_l1_done;
        prev_goodness_l2_done <= dut.goodness_l2_done;

        // Detect rising edge of goodness_l2_done
        if (dut.goodness_l2_done && !prev_goodness_l2_done) begin
            if (dut.ctrl.fwd_state == 8) begin  // FWD_L2_GOODNESS
                if (dut.ctrl.is_positive_pass) begin
                    pos_goodness_f = q_to_real(dut.goodness_l2_val);
                    $fdisplay(log_file, "%0d,pos,%.4f",
                              sample_count, pos_goodness_f);
                end
                else begin
                    neg_goodness_f = q_to_real(dut.goodness_l2_val);
                    $fdisplay(log_file, "%0d,neg,%.4f",
                              sample_count, neg_goodness_f);
                    // Both passes done for this sample — print summary
                    $display("[TB] Sample %4d | Pos: %7.3f | Neg: %7.3f",
                             sample_count,
                             q_to_real(dut.goodness_l2_val),
                             neg_goodness_f);
                    sample_count <= sample_count + 1;
                end
            end
        end
    end

    // ─────────────────────────────────────────────
    // WEIGHT CHANGE MONITOR
    // Verify learning is happening by checking
    // that weights are actually changing
    // Samples spot-check weights at fixed addresses
    // ─────────────────────────────────────────────
    logic [DATA_WIDTH-1:0] w1_spot_before;
    logic [DATA_WIDTH-1:0] w2_spot_before;
    localparam SPOT_ADDR_L1 = 100;   // arbitrary weight addresses to watch
    localparam SPOT_ADDR_L2 = 50;

    task capture_spot_weights();
        w1_spot_before = dut.l1_wbram.mem[SPOT_ADDR_L1];
        w2_spot_before = dut.l2_wbram.mem[SPOT_ADDR_L2];
        $display("[TB] Spot weights before training:");
        $display("     L1[%0d] = %h (%.4f)",
                 SPOT_ADDR_L1, w1_spot_before,
                 q_to_real(w1_spot_before));
        $display("     L2[%0d] = %h (%.4f)",
                 SPOT_ADDR_L2, w2_spot_before,
                 q_to_real(w2_spot_before));
    endtask

    task check_spot_weights();
        logic [DATA_WIDTH-1:0] w1_after, w2_after;
        w1_after = dut.l1_wbram.mem[SPOT_ADDR_L1];
        w2_after = dut.l2_wbram.mem[SPOT_ADDR_L2];
        $display("[TB] Spot weights after training:");
        $display("     L1[%0d] = %h (%.4f)",
                 SPOT_ADDR_L1, w1_after,
                 q_to_real(w1_after));
        $display("     L2[%0d] = %h (%.4f)",
                 SPOT_ADDR_L2, w2_after,
                 q_to_real(w2_after));

        if (w1_after !== w1_spot_before)
            $display("[TB] PASS: L1 weights changed — learning confirmed.");
        else
            $display("[TB] FAIL: L1 weights unchanged — learning not happening.");

        if (w2_after !== w2_spot_before)
            $display("[TB] PASS: L2 weights changed — learning confirmed.");
        else
            $display("[TB] FAIL: L2 weights unchanged — learning not happening.");
    endtask

    // ─────────────────────────────────────────────
    // SAMPLE MEMORY LOADER
    // Converts Python mem_files format to
    // flat sample_mem array
    // Python exports one sample per row of 784 values
    // Testbench expects flat: sample 0 pixel 0..783,
    // then sample 1 pixel 0..783, etc.
    // ─────────────────────────────────────────────
    task load_samples();
        $display("[TB] Loading MNIST samples from mem_files/...");
        // Load first NUM_SAMPLES images from full dataset mem file
        // Python should export samples_flat.mem with all pixels
        // in row-major order: s0p0, s0p1...s0p783, s1p0...
        $readmemh("C:/Users/youss/Documents/Forward-Forward-RTL-Implementation-w-Parallel-Inference-and-Training/mem_files/samples_flat.mem", sample_mem, 0, (NUM_SAMPLES * L1_INPUT_SIZE) - 1);
        $readmemh("C:/Users/youss/Documents/Forward-Forward-RTL-Implementation-w-Parallel-Inference-and-Training/mem_files/labels.mem", label_mem, 0, NUM_SAMPLES - 1);
        $display("[TB] Samples loaded.");
        $display("[TB] Samples loaded.");
    endtask

    // ─────────────────────────────────────────────
    // PARALLEL DATAPATH MONITOR
    // Verifies the key architectural claim:
    // PE_L1 and L2_MAC actually overlap in time.
    // Records timestamps when each starts and ends.
    // ─────────────────────────────────────────────
    longint pe_l1_start_time,  pe_l1_end_time;
    longint l2_mac_start_time, l2_mac_end_time;
    logic   pe_l1_started, l2_mac_started;
    logic   overlap_confirmed;

    always_ff @(posedge clk) begin
        // Detect PE starting on layer 1
        if (dut.pe_start && !dut.pe_layer_sel && !pe_l1_started) begin
            pe_l1_start_time <= $time;
            pe_l1_started    <= 1'b1;
        end
        if (dut.pe_done && pe_l1_started && !dut.pe_layer_sel) begin
            pe_l1_end_time <= $time;
            pe_l1_started  <= 1'b0;
        end

        // Detect L2 MAC starting
        if (dut.l2_mac_start && !l2_mac_started) begin
            l2_mac_start_time <= $time;
            l2_mac_started    <= 1'b1;
        end
        if (dut.l2_mac_done && l2_mac_started) begin
            l2_mac_end_time <= $time;
            l2_mac_started  <= 1'b0;

            // Check overlap: L2 MAC started before PE_L1 ended
            if (l2_mac_start_time >= pe_l1_start_time &&
                l2_mac_start_time <= pe_l1_end_time) begin
                if (!overlap_confirmed) begin
                    $display("[TB] PARALLEL CONFIRMED: L2_MAC started at %0t",
                             l2_mac_start_time);
                    $display("     PE_L1 was running from %0t to %0t",
                             pe_l1_start_time, pe_l1_end_time);
                    $display("     Overlap = %0t ns",
                             pe_l1_end_time - l2_mac_start_time);
                    overlap_confirmed <= 1'b1;
                end
            end
        end
    end

    // ─────────────────────────────────────────────
    // MAIN STIMULUS
    // ─────────────────────────────────────────────
    integer chk;

    initial begin
        // ── SETUP ─────────────────────────────────
        $display("================================================");
        $display("  Forward-Forward RTL Testbench");
        $display("  Architecture: 784->256->256");
        $display("  Samples: %0d", NUM_SAMPLES);
        $display("  Clock: 100MHz");
        $display("================================================");

        // Open log file for goodness tracking
        log_file = $fopen("sim_goodness_log.csv", "w");
        $fdisplay(log_file, "sample,pass,goodness");

        // Initialize tracking variables
        checkpoint_num  <= 0;
        in_positive_pass  <= 1'b1;

        // Initialize signals
        rst_n = 0;
        start = 0;

        // ── RESET ─────────────────────────────────
        repeat(10) @(posedge clk);
        rst_n = 1;
        repeat(5) @(posedge clk);

        // ── LOAD MEMORIES ─────────────────────────
        load_samples();
        load_weights();
        capture_spot_weights();

        // Create checkpoints directory
        // Note: $system may not work in all simulators
        // Create manually if needed
        $display("[TB] Starting training...");
        repeat(5) @(posedge clk);

        // ── START TRAINING ────────────────────────
        @(posedge clk);
        start = 1;
        @(posedge clk);
        start = 0;

        // ── WAIT FOR COMPLETION ───────────────────
        // Poll for training_done with timeout
        // Timeout = 2B cycles at 100MHz = 20 seconds sim time
        fork
            begin : wait_done
                wait(training_done);
                $display("[TB] training_done received at time %0t", $time);
                disable timeout_block;
            end
            begin : timeout_block
                repeat(2_000_000_000) @(posedge clk);
                $display("[TB] TIMEOUT — training did not complete.");
                disable wait_done;
            end
        join

        // ── POST-TRAINING CHECKS ──────────────────
        repeat(10) @(posedge clk);

        $display("");
        $display("================================================");
        $display("  Training Complete — Results");
        $display("================================================");

        // Verify weights changed
        check_spot_weights();

        // Final weight dump
        dump_weights(99);

        // Report parallel overlap
        if (overlap_confirmed)
            $display("[TB] Dual-datapath parallelism: VERIFIED");
        else
            $display("[TB] Dual-datapath parallelism: NOT OBSERVED — check FSM");

        // Close log
        $fclose(log_file);

        $display("");
        $display("[TB] Goodness log written to sim_goodness_log.csv");
        $display("[TB] Final weights written to checkpoints/chk99_layer*.mem");
        $display("[TB] Done.");
        $display("================================================");

        $finish;
    end

    // ─────────────────────────────────────────────
    // PERIODIC CHECKPOINT TASK
    // Triggered by sample_count advancing
    // ─────────────────────────────────────────────
    always_ff @(posedge clk) begin
        if (sample_count > 0 &&
            sample_count % CHECKPOINT_INTERVAL == 0 &&
            !dut.ctrl.is_positive_pass) begin
            dump_weights(sample_count / CHECKPOINT_INTERVAL);
        end
    end

    // ─────────────────────────────────────────────
    // WAVEFORM DUMP
    // Captures key signals for ModelSim waveform view
    // Add signals you want to watch here
    // ─────────────────────────────────────────────
    initial begin
        $dumpfile("ff_sim.vcd");
        $dumpvars(0, tb_top);
    end

endmodule
